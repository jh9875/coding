-- week10_class2.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY week10_class2 IS
PORT(
	RESETN : IN STD_LOGIC;
	CLK : IN STD_LOGIC;
	
    BCD : IN STD_LOGIC_VECTOR(15 downto 0);
    a, b, c, d, e, f, g : OUT STD_LOGIC;
	PIEZO : OUT STD_LOGIC
);
END week10_class2;

ARCHITECTURE HB OF week10_class2 IS

	SIGNAL DECODE : STD_LOGIC_VECTOR(6 downto 0);
	
	CONSTANT CNT_DO : INTEGER RANGE 0 TO 2047 := 1910;     
	CONSTANT CNT_RAE : INTEGER RANGE 0 TO 2047 := 1701;      
	CONSTANT CNT_MI : INTEGER RANGE 0 TO 2047 := 1516;     
	CONSTANT CNT_FA : INTEGER RANGE 0 TO 2047 := 1431;     
	CONSTANT CNT_SOL : INTEGER RANGE 0 TO 2047 := 1275;     
	CONSTANT CNT_RA : INTEGER RANGE 0 TO 2047 := 1135;     
	CONSTANT CNT_SI : INTEGER RANGE 0 TO 2047 := 1011;     
	CONSTANT CNT_HDO : INTEGER RANGE 0 TO 2047 := 955; 
 
	SIGNAL REG : STD_LOGIC;
	SIGNAL CNT : INTEGER RANGE 0 TO 2047;     
	SIGNAL LIMIT : INTEGER RANGE 0 TO 2047; 

BEGIN

-- 버튼에 해당하는 음계의 소리를 내도록 지정
PROCESS(BCD) 
BEGIN     
	CASE BCD IS    -- 이 부분도 수정
		WHEN "0000000000000001" => LIMIT <= 1910;    -- 도
		WHEN "0000000000000010" => LIMIT <= 1701;    -- 레
		WHEN "0000000000000100" => LIMIT <= 1516;    -- 미
		WHEN "0000000000001000" => LIMIT <= 1431;   -- 파
		WHEN "0000000000010000" => LIMIT <= 1275;    -- 솔
		WHEN "0000000000100000" => LIMIT <= 1135;     -- 라
		WHEN "0000000001000000" => LIMIT <= 1011;    -- 시
		WHEN "0000000010000000" => LIMIT <= 955;    -- 높은 도
		WHEN OTHERS => LIMIT <= 0;  
	END CASE; 
END PROCESS; 

-- 클럭이 발생하였을 때, 
-- 주파수 생성을 위한 카운트 하는 변수 CNT를 앞에서 설정한 LIMIT까지 카운트하여 
-- REG 주파수를 생성
-- 이 코드는 건들일 필요 없음.
PROCESS(RESETN, CLK) 
BEGIN  
   IF RESETN = '0' THEN 
	    CNT <= 0;     
	    REG <= '0';   
   ELSIF CLK'EVENT AND CLK = '1' THEN  
		IF CNT >= LIMIT THEN           
			CNT <= 0;         
			REG <= NOT REG;     
	    ELSE           
			CNT <= CNT + 1;      
	    END IF;  
   END IF; 
END PROCESS; 
 
-- 세그먼트 PROCESS

PROCESS(BCD)
BEGIN
    CASE BCD IS
        WHEN "0000001000000000" => DECODE <= "1111110";
        WHEN "0000000000000001" => DECODE <= "0110000"; -- 1
        WHEN "0000000000000010" => DECODE <= "1101101"; -- 2
        WHEN "0000000000000100" => DECODE <= "1111001"; -- 3
        WHEN "0000000000001000" => DECODE <= "0110011"; -- 4
        WHEN "0000000000010000" => DECODE <= "1011011"; -- 5
        WHEN "0000000000100000" => DECODE <= "1011111"; -- 6
        WHEN "0000000001000000" => DECODE <= "1110000"; -- 7
        WHEN "0000000010000000" => DECODE <= "1111111"; -- 8
        WHEN "0000000100000000" => DECODE <= "1111011"; -- 9
        WHEN "0000010000000000" => DECODE <= "1110111"; -- A
	    WHEN "0000100000000000" => DECODE <= "0011111"; -- B
	    WHEN "0001000000000000" => DECODE <= "1001110"; -- C
	    WHEN "0010000000000000" => DECODE <= "0111101"; -- D
	    WHEN "0100000000000000" => DECODE <= "1001111"; -- E
	    WHEN "1000000000000000" => DECODE <= "1000111"; -- F		  
        WHEN OTHERS => NULL;
    END CASE;
END PROCESS;

a <= DECODE(6);
b <= DECODE(5);
c <= DECODE(4);
d <= DECODE(3);
e <= DECODE(2);
f <= DECODE(1);
g <= DECODE(0);

PIEZO <= REG;
 

END HB;