-- HB_SEG_DISP.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY HB_SEG_DISP IS
	PORT(
		RESETN   : IN  STD_LOGIC;       -- RESET
		CLK      : IN  STD_LOGIC;       -- 1kHz CLOCK
		SEG_COM  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- 7-SEGMENT COMMON SELECT
		SEG_DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) -- 7-SEGMENT DATA
	);
END HB_SEG_DISP;

ARCHITECTURE HB OF HB_SEG_DISP IS
	SIGNAL CNT_SCAN : INTEGER RANGE 0 TO 3; -- SCAN COUNT

BEGIN
	-- SCAN COUNT
	PROCESS(RESETN, CLK)
	BEGIN
		IF RESETN = '0' THEN
			CNT_SCAN <= 0;
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF CNT_SCAN = 3 THEN
				CNT_SCAN <= 0;
			ELSE
				CNT_SCAN <= CNT_SCAN + 1;
			END IF;
		END IF;
	END PROCESS;

	-- SEGMENT DISPLAY
	PROCESS(RESETN, CLK)
	BEGIN
		IF RESETN = '0' THEN
			SEG_COM  <= X"FF";
			SEG_DATA <= X"00";
		ELSIF CLK'EVENT AND CLK = '1' THEN
			CASE CNT_SCAN IS
				WHEN 0 =>
					SEG_COM  <= X"7";   -- SEL COM1
					SEG_DATA <= X"C";   -- 0
				WHEN 1 =>
					SEG_COM  <= X"B";   -- SEL COM2
					SEG_DATA <= X"60";  -- 1
				WHEN 2 =>
					SEG_COM  <= X"D";   -- SEL COM3
					SEG_DATA <= X"DA";  -- 2
				WHEN 3 =>
					SEG_COM  <= X"E";   -- SEL COM4
					SEG_DATA <= X"F2";  -- 3
				WHEN OTHERS =>
					SEG_COM  <= X"F";   -- SEL X
					SEG_DATA <= X"00";  --
			END CASE;
		END IF;
	END PROCESS;
END HB;
