--TB_HB_OR2.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_XNOR IS
END TB_HB_XNOR;

ARCHITECTURE HB OF TB_HB_XNOR IS
	COMPONENT HB_XNOR
		PORT(
			A, B, C : IN  BIT;
			X    : OUT BIT
		);
	END COMPONENT;
	SIGNAL A : BIT := '0';
	SIGNAL B : BIT := '0';
	SIGNAL C : BIT := '0';
	SIGNAL X : BIT := '0';
BEGIN
	A <= '0', '1' AFTER 400 NS;
	B <= '0', '1' AFTER 200 NS, '0' AFTER 400 NS, '1' AFTER 600 NS;
	C <= '0', '1' AFTER 100 NS, '0' AFTER 200 NS, '1' AFTER 300 NS, '0' AFTER 400 NS, '1' AFTER 500 NS, '0' AFTER 600 NS,
			'1' AFTER 700 NS, '0' AFTER 800 NS;
	U_HB_XNOR : HB_XNOR
		PORT MAP(
			A => A,
			B => B,
			C => C,
			X => X
		);
END HB;
