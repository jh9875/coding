--TB_HB_HS.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_HS IS
END TB_HB_HS;

ARCHITECTURE HB OF TB_HB_HS IS
	COMPONENT HB_HS
		PORT(
			A, B : IN  BIT;
			D, B0 : OUT BIT
		);
	END COMPONENT;

	SIGNAL A, B : BIT := '0';
	SIGNAL D, B0 : BIT := '0';

BEGIN
	A <= '0', '1' AFTER 200 NS;
	B <= '0', '1' AFTER 100 NS, '0' AFTER 200 NS, '1' AFTER 300 NS, '0' AFTER 400 NS;
	U_HB_HS : HB_HS
		PORT MAP(
			A => A,
			B => B,
			D => D,
			B0 => B0
		);
END HB;
